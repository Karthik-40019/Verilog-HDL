`timescale 1ns/100ps

module cmos_fullAdder_tb;
reg a,b,cin;
wire sum,cout;

cmos_fullAdder uut(a,b,cin,sum,cout);
initial begin 

a=0;b=0;cin=0;#10;
a=0;b=0;cin=1;#10;
a=0;b=1;cin=0;#10;
a=0;b=1;cin=1;#10;

a=1;b=0;cin=0;#10;
a=1;b=0;cin=1;#10;
a=1;b=1;cin=0;#10;
a=1;b=1;cin=1;#10;

end
endmodule
